`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/13 19:36:20
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module top(
input clk,
input rst,
input [6:0] fp7_0_A0,input [6:0] fp7_0_B0,
input [6:0] fp7_0_A1,input [6:0] fp7_0_B1,
input [6:0] fp7_0_A2,input [6:0] fp7_0_B2,
input [6:0] fp7_0_A3,input [6:0] fp7_0_B3,
input [6:0] fp7_0_A4,input [6:0] fp7_0_B4,
input [6:0] fp7_0_A5,input [6:0] fp7_0_B5,
input [6:0] fp7_0_A6,input [6:0] fp7_0_B6,
input [6:0] fp7_0_A7,input [6:0] fp7_0_B7,
input [1:0]fp7_0_sig0,input [1:0]fp7_0_sig1,
input [1:0]fp7_0_sig2,input [1:0]fp7_0_sig3,
input [1:0]fp7_0_sig4,input [1:0]fp7_0_sig5,
input [1:0]fp7_0_sig6,input [1:0]fp7_0_sig7,
input [7:0]fp7_0_exp0,input [7:0]fp7_0_exp1,
input [7:0]fp7_0_exp2,input [7:0]fp7_0_exp3,
input [7:0]fp7_0_exp4,input [7:0]fp7_0_exp5,
input [7:0]fp7_0_exp6,input [7:0]fp7_0_exp7,
output [31:0] fp7_0_out,

input [6:0] fp7_1_A0,input [6:0] fp7_1_B0,
input [6:0] fp7_1_A1,input [6:0] fp7_1_B1,
input [6:0] fp7_1_A2,input [6:0] fp7_1_B2,
input [6:0] fp7_1_A3,input [6:0] fp7_1_B3,
input [6:0] fp7_1_A4,input [6:0] fp7_1_B4,
input [6:0] fp7_1_A5,input [6:0] fp7_1_B5,
input [6:0] fp7_1_A6,input [6:0] fp7_1_B6,
input [6:0] fp7_1_A7,input [6:0] fp7_1_B7,
input [1:0]fp7_1_sig0,input [1:0]fp7_1_sig1,
input [1:0]fp7_1_sig2,input [1:0]fp7_1_sig3,
input [1:0]fp7_1_sig4,input [1:0]fp7_1_sig5,
input [1:0]fp7_1_sig6,input [1:0]fp7_1_sig7,
input [7:0]fp7_1_exp0,input [7:0]fp7_1_exp1,
input [7:0]fp7_1_exp2,input [7:0]fp7_1_exp3,
input [7:0]fp7_1_exp4,input [7:0]fp7_1_exp5,
input [7:0]fp7_1_exp6,input [7:0]fp7_1_exp7,
output [31:0] fp7_1_out,

input [6:0] fp7_2_A0,input [6:0] fp7_2_B0,
input [6:0] fp7_2_A1,input [6:0] fp7_2_B1,
input [6:0] fp7_2_A2,input [6:0] fp7_2_B2,
input [6:0] fp7_2_A3,input [6:0] fp7_2_B3,
input [6:0] fp7_2_A4,input [6:0] fp7_2_B4,
input [6:0] fp7_2_A5,input [6:0] fp7_2_B5,
input [6:0] fp7_2_A6,input [6:0] fp7_2_B6,
input [6:0] fp7_2_A7,input [6:0] fp7_2_B7,
input [1:0]fp7_2_sig0,input [1:0]fp7_2_sig1,
input [1:0]fp7_2_sig2,input [1:0]fp7_2_sig3,
input [1:0]fp7_2_sig4,input [1:0]fp7_2_sig5,
input [1:0]fp7_2_sig6,input [1:0]fp7_2_sig7,
input [7:0]fp7_2_exp0,input [7:0]fp7_2_exp1,
input [7:0]fp7_2_exp2,input [7:0]fp7_2_exp3,
input [7:0]fp7_2_exp4,input [7:0]fp7_2_exp5,
input [7:0]fp7_2_exp6,input [7:0]fp7_2_exp7,
output [31:0] fp7_2_out,

input [8:0] fp8_0_A0,input [8:0] fp8_0_B0,
input [8:0] fp8_0_A1,input [8:0] fp8_0_B1,
input [8:0] fp8_0_A2,input [8:0] fp8_0_B2,
input [8:0] fp8_0_A3,input [8:0] fp8_0_B3,
input [8:0] fp8_0_A4,input [8:0] fp8_0_B4,
input [8:0] fp8_0_A5,input [8:0] fp8_0_B5,
input [8:0] fp8_0_A6,input [8:0] fp8_0_B6,
input [8:0] fp8_0_A7,input [8:0] fp8_0_B7,
output [31:0] fp8_0_out,

input [8:0] fp8_1_A0,input [8:0] fp8_1_B0,
input [8:0] fp8_1_A1,input [8:0] fp8_1_B1,
input [8:0] fp8_1_A2,input [8:0] fp8_1_B2,
input [8:0] fp8_1_A3,input [8:0] fp8_1_B3,
input [8:0] fp8_1_A4,input [8:0] fp8_1_B4,
input [8:0] fp8_1_A5,input [8:0] fp8_1_B5,
input [8:0] fp8_1_A6,input [8:0] fp8_1_B6,
input [8:0] fp8_1_A7,input [8:0] fp8_1_B7,
output [31:0] fp8_1_out,

input [8:0] fp8_2_A0,input [8:0] fp8_2_B0,
input [8:0] fp8_2_A1,input [8:0] fp8_2_B1,
input [8:0] fp8_2_A2,input [8:0] fp8_2_B2,
input [8:0] fp8_2_A3,input [8:0] fp8_2_B3,
input [8:0] fp8_2_A4,input [8:0] fp8_2_B4,
input [8:0] fp8_2_A5,input [8:0] fp8_2_B5,
input [8:0] fp8_2_A6,input [8:0] fp8_2_B6,
input [8:0] fp8_2_A7,input [8:0] fp8_2_B7,
output [31:0] fp8_2_out,

input [31:0] fp32_0_A0,input [31:0] fp32_0_B0,
input [31:0] fp32_0_A1,input [31:0] fp32_0_B1,
input [31:0] fp32_0_A2,input [31:0] fp32_0_B2,
input [31:0] fp32_0_A3,input [31:0] fp32_0_B3,
input [31:0] fp32_0_A4,input [31:0] fp32_0_B4,
input [31:0] fp32_0_A5,input [31:0] fp32_0_B5,
input [31:0] fp32_0_A6,input [31:0] fp32_0_B6,
input [31:0] fp32_0_A7,input [31:0] fp32_0_B7,
output [31:0] fp32_0_out,

input [31:0] fp32_1_A0,input [31:0] fp32_1_B0,
input [31:0] fp32_1_A1,input [31:0] fp32_1_B1,
input [31:0] fp32_1_A2,input [31:0] fp32_1_B2,
input [31:0] fp32_1_A3,input [31:0] fp32_1_B3,
input [31:0] fp32_1_A4,input [31:0] fp32_1_B4,
input [31:0] fp32_1_A5,input [31:0] fp32_1_B5,
input [31:0] fp32_1_A6,input [31:0] fp32_1_B6,
input [31:0] fp32_1_A7,input [31:0] fp32_1_B7,
output [31:0] fp32_1_out,

input [31:0] fp32_2_A0,input [31:0] fp32_2_B0,
input [31:0] fp32_2_A1,input [31:0] fp32_2_B1,
input [31:0] fp32_2_A2,input [31:0] fp32_2_B2,
input [31:0] fp32_2_A3,input [31:0] fp32_2_B3,
input [31:0] fp32_2_A4,input [31:0] fp32_2_B4,
input [31:0] fp32_2_A5,input [31:0] fp32_2_B5,
input [31:0] fp32_2_A6,input [31:0] fp32_2_B6,
input [31:0] fp32_2_A7,input [31:0] fp32_2_B7,
output [31:0] fp32_2_out,

input [7:0] int8_0_A0,input [7:0] int8_0_B0,
input [7:0] int8_0_A1,input [7:0] int8_0_B1,
input [7:0] int8_0_A2,input [7:0] int8_0_B2,
input [7:0] int8_0_A3,input [7:0] int8_0_B3,
input [7:0] int8_0_A4,input [7:0] int8_0_B4,
input [7:0] int8_0_A5,input [7:0] int8_0_B5,
input [7:0] int8_0_A6,input [7:0] int8_0_B6,
input [7:0] int8_0_A7,input [7:0] int8_0_B7,
output [31:0] int8_0_out,

input [7:0] int8_1_A0,input [7:0] int8_1_B0,
input [7:0] int8_1_A1,input [7:0] int8_1_B1,
input [7:0] int8_1_A2,input [7:0] int8_1_B2,
input [7:0] int8_1_A3,input [7:0] int8_1_B3,
input [7:0] int8_1_A4,input [7:0] int8_1_B4,
input [7:0] int8_1_A5,input [7:0] int8_1_B5,
input [7:0] int8_1_A6,input [7:0] int8_1_B6,
input [7:0] int8_1_A7,input [7:0] int8_1_B7,
output [31:0] int8_1_out,

input [7:0] int8_2_A0,input [7:0] int8_2_B0,
input [7:0] int8_2_A1,input [7:0] int8_2_B1,
input [7:0] int8_2_A2,input [7:0] int8_2_B2,
input [7:0] int8_2_A3,input [7:0] int8_2_B3,
input [7:0] int8_2_A4,input [7:0] int8_2_B4,
input [7:0] int8_2_A5,input [7:0] int8_2_B5,
input [7:0] int8_2_A6,input [7:0] int8_2_B6,
input [7:0] int8_2_A7,input [7:0] int8_2_B7,
output [31:0] int8_2_out,

input [1:0] mulPE_0_ctrl,
input [31:0] mulPE_0_scalar,
input [31:0] mulPE_0_A0,input [31:0] mulPE_0_B0,
input [31:0] mulPE_0_A1,input [31:0] mulPE_0_B1,
input [31:0] mulPE_0_A2,input [31:0] mulPE_0_B2,
input [31:0] mulPE_0_A3,input [31:0] mulPE_0_B3,
input [31:0] mulPE_0_A4,input [31:0] mulPE_0_B4,
input [31:0] mulPE_0_A5,input [31:0] mulPE_0_B5,
input [31:0] mulPE_0_A6,input [31:0] mulPE_0_B6,
input [31:0] mulPE_0_A7,input [31:0] mulPE_0_B7,
output [31:0] mulPE_0_out0,
output [31:0] mulPE_0_out1,
output [31:0] mulPE_0_out2,
output [31:0] mulPE_0_out3,
output [31:0] mulPE_0_out4,
output [31:0] mulPE_0_out5,
output [31:0] mulPE_0_out6,
output [31:0] mulPE_0_out7,

input [1:0] mulPE_1_ctrl,
input [31:0] mulPE_1_scalar,
input [31:0] mulPE_1_A0,input [31:0] mulPE_1_B0,
input [31:0] mulPE_1_A1,input [31:0] mulPE_1_B1,
input [31:0] mulPE_1_A2,input [31:0] mulPE_1_B2,
input [31:0] mulPE_1_A3,input [31:0] mulPE_1_B3,
input [31:0] mulPE_1_A4,input [31:0] mulPE_1_B4,
input [31:0] mulPE_1_A5,input [31:0] mulPE_1_B5,
input [31:0] mulPE_1_A6,input [31:0] mulPE_1_B6,
input [31:0] mulPE_1_A7,input [31:0] mulPE_1_B7,
output [31:0] mulPE_1_out0,
output [31:0] mulPE_1_out1,
output [31:0] mulPE_1_out2,
output [31:0] mulPE_1_out3,
output [31:0] mulPE_1_out4,
output [31:0] mulPE_1_out5,
output [31:0] mulPE_1_out6,
output [31:0] mulPE_1_out7,

input [1:0] mulPE_2_ctrl,
input [31:0] mulPE_2_scalar,
input [31:0] mulPE_2_A0,input [31:0] mulPE_2_B0,
input [31:0] mulPE_2_A1,input [31:0] mulPE_2_B1,
input [31:0] mulPE_2_A2,input [31:0] mulPE_2_B2,
input [31:0] mulPE_2_A3,input [31:0] mulPE_2_B3,
input [31:0] mulPE_2_A4,input [31:0] mulPE_2_B4,
input [31:0] mulPE_2_A5,input [31:0] mulPE_2_B5,
input [31:0] mulPE_2_A6,input [31:0] mulPE_2_B6,
input [31:0] mulPE_2_A7,input [31:0] mulPE_2_B7,
output [31:0] mulPE_2_out0,
output [31:0] mulPE_2_out1,
output [31:0] mulPE_2_out2,
output [31:0] mulPE_2_out3,
output [31:0] mulPE_2_out4,
output [31:0] mulPE_2_out5,
output [31:0] mulPE_2_out6,
output [31:0] mulPE_2_out7,

input addPE_0_ctrl,
input [31:0] addPE_0_scalar,
input [31:0] addPE_0_A0,input [31:0] addPE_0_B0,
input [31:0] addPE_0_A1,input [31:0] addPE_0_B1,
input [31:0] addPE_0_A2,input [31:0] addPE_0_B2,
input [31:0] addPE_0_A3,input [31:0] addPE_0_B3,
input [31:0] addPE_0_A4,input [31:0] addPE_0_B4,
input [31:0] addPE_0_A5,input [31:0] addPE_0_B5,
input [31:0] addPE_0_A6,input [31:0] addPE_0_B6,
input [31:0] addPE_0_A7,input [31:0] addPE_0_B7,
output [31:0] addPE_0_out0,
output [31:0] addPE_0_out1,
output [31:0] addPE_0_out2,
output [31:0] addPE_0_out3,
output [31:0] addPE_0_out4,
output [31:0] addPE_0_out5,
output [31:0] addPE_0_out6,
output [31:0] addPE_0_out7,

input addPE_1_ctrl,
input [31:0] addPE_1_scalar,
input [31:0] addPE_1_A0,input [31:0] addPE_1_B0,
input [31:0] addPE_1_A1,input [31:0] addPE_1_B1,
input [31:0] addPE_1_A2,input [31:0] addPE_1_B2,
input [31:0] addPE_1_A3,input [31:0] addPE_1_B3,
input [31:0] addPE_1_A4,input [31:0] addPE_1_B4,
input [31:0] addPE_1_A5,input [31:0] addPE_1_B5,
input [31:0] addPE_1_A6,input [31:0] addPE_1_B6,
input [31:0] addPE_1_A7,input [31:0] addPE_1_B7,
output [31:0] addPE_1_out0,
output [31:0] addPE_1_out1,
output [31:0] addPE_1_out2,
output [31:0] addPE_1_out3,
output [31:0] addPE_1_out4,
output [31:0] addPE_1_out5,
output [31:0] addPE_1_out6,
output [31:0] addPE_1_out7,

input addPE_2_ctrl,
input [31:0] addPE_2_scalar,
input [31:0] addPE_2_A0,input [31:0] addPE_2_B0,
input [31:0] addPE_2_A1,input [31:0] addPE_2_B1,
input [31:0] addPE_2_A2,input [31:0] addPE_2_B2,
input [31:0] addPE_2_A3,input [31:0] addPE_2_B3,
input [31:0] addPE_2_A4,input [31:0] addPE_2_B4,
input [31:0] addPE_2_A5,input [31:0] addPE_2_B5,
input [31:0] addPE_2_A6,input [31:0] addPE_2_B6,
input [31:0] addPE_2_A7,input [31:0] addPE_2_B7,
output [31:0] addPE_2_out0,
output [31:0] addPE_2_out1,
output [31:0] addPE_2_out2,
output [31:0] addPE_2_out3,
output [31:0] addPE_2_out4,
output [31:0] addPE_2_out5,
output [31:0] addPE_2_out6,
output [31:0] addPE_2_out7,

input [31:0] treePE_0_A0,
input [31:0] treePE_0_A1,
input [31:0] treePE_0_A2,
input [31:0] treePE_0_A3,
input [31:0] treePE_0_A4,
input [31:0] treePE_0_A5,
input [31:0] treePE_0_A6,
input [31:0] treePE_0_A7,
output[31:0] treePE_0_out,

input [31:0] treePE_1_A0,
input [31:0] treePE_1_A1,
input [31:0] treePE_1_A2,
input [31:0] treePE_1_A3,
input [31:0] treePE_1_A4,
input [31:0] treePE_1_A5,
input [31:0] treePE_1_A6,
input [31:0] treePE_1_A7,
output[31:0] treePE_1_out,

input [31:0] treePE_2_A0,
input [31:0] treePE_2_A1,
input [31:0] treePE_2_A2,
input [31:0] treePE_2_A3,
input [31:0] treePE_2_A4,
input [31:0] treePE_2_A5,
input [31:0] treePE_2_A6,
input [31:0] treePE_2_A7,
output[31:0] treePE_2_out



);

fp7PE fp7_0(
    clk,rst,
fp7_0_A0,fp7_0_B0,
fp7_0_A1,fp7_0_B1,
fp7_0_A2,fp7_0_B2,
fp7_0_A3,fp7_0_B3,
fp7_0_A4,fp7_0_B4,
fp7_0_A5,fp7_0_B5,
fp7_0_A6,fp7_0_B6,
fp7_0_A7,fp7_0_B7,
fp7_0_sig0,fp7_0_sig1,
fp7_0_sig2,fp7_0_sig3,
fp7_0_sig4,fp7_0_sig5,
fp7_0_sig6,fp7_0_sig7,
fp7_0_exp0,fp7_0_exp1,
fp7_0_exp2,fp7_0_exp3,
fp7_0_exp4,fp7_0_exp5,
fp7_0_exp6,fp7_0_exp7,
fp7_0_out);

fp7PE fp7_1(
    clk,rst,
fp7_1_A0,fp7_1_B0,
fp7_1_A1,fp7_1_B1,
fp7_1_A2,fp7_1_B2,
fp7_1_A3,fp7_1_B3,
fp7_1_A4,fp7_1_B4,
fp7_1_A5,fp7_1_B5,
fp7_1_A6,fp7_1_B6,
fp7_1_A7,fp7_1_B7,
fp7_1_sig0,fp7_1_sig1,
fp7_1_sig2,fp7_1_sig3,
fp7_1_sig4,fp7_1_sig5,
fp7_1_sig6,fp7_1_sig7,
fp7_1_exp0,fp7_1_exp1,
fp7_1_exp2,fp7_1_exp3,
fp7_1_exp4,fp7_1_exp5,
fp7_1_exp6,fp7_1_exp7,
fp7_1_out);

fp7PE fp7_2(clk,rst,
fp7_2_A0,fp7_2_B0,
fp7_2_A1,fp7_2_B1,
fp7_2_A2,fp7_2_B2,
fp7_2_A3,fp7_2_B3,
fp7_2_A4,fp7_2_B4,
fp7_2_A5,fp7_2_B5,
fp7_2_A6,fp7_2_B6,
fp7_2_A7,fp7_2_B7,
fp7_2_sig0,fp7_2_sig1,
fp7_2_sig2,fp7_2_sig3,
fp7_2_sig4,fp7_2_sig5,
fp7_2_sig6,fp7_2_sig7,
fp7_2_exp0,fp7_2_exp1,
fp7_2_exp2,fp7_2_exp3,
fp7_2_exp4,fp7_2_exp5,
fp7_2_exp6,fp7_2_exp7,
fp7_2_out);

fp8PE fp8_0(clk,rst,
fp8_0_A0,fp8_0_B0,
fp8_0_A1,fp8_0_B1,
fp8_0_A2,fp8_0_B2,
fp8_0_A3,fp8_0_B3,
fp8_0_A4,fp8_0_B4,
fp8_0_A5,fp8_0_B5,
fp8_0_A6,fp8_0_B6,
fp8_0_A7,fp8_0_B7,
fp8_0_out
);

fp8PE fp8_1(clk,rst,
fp8_1_A0,fp8_1_B0,
fp8_1_A1,fp8_1_B1,
fp8_1_A2,fp8_1_B2,
fp8_1_A3,fp8_1_B3,
fp8_1_A4,fp8_1_B4,
fp8_1_A5,fp8_1_B5,
fp8_1_A6,fp8_1_B6,
fp8_1_A7,fp8_1_B7,
fp8_1_out
);

fp8PE fp8_2(clk,rst,
fp8_2_A0,fp8_2_B0,
fp8_2_A1,fp8_2_B1,
fp8_2_A2,fp8_2_B2,
fp8_2_A3,fp8_2_B3,
fp8_2_A4,fp8_2_B4,
fp8_2_A5,fp8_2_B5,
fp8_2_A6,fp8_2_B6,
fp8_2_A7,fp8_2_B7,
fp8_2_out
);

fp32PE fp32_0(clk,rst,
fp32_0_A0,fp32_0_B0,
fp32_0_A1,fp32_0_B1,
fp32_0_A2,fp32_0_B2,
fp32_0_A3,fp32_0_B3,
fp32_0_A4,fp32_0_B4,
fp32_0_A5,fp32_0_B5,
fp32_0_A6,fp32_0_B6,
fp32_0_A7,fp32_0_B7,
fp32_0_out
);

fp32PE fp32_1(clk,rst,
fp32_1_A0,fp32_1_B0,
fp32_1_A1,fp32_1_B1,
fp32_1_A2,fp32_1_B2,
fp32_1_A3,fp32_1_B3,
fp32_1_A4,fp32_1_B4,
fp32_1_A5,fp32_1_B5,
fp32_1_A6,fp32_1_B6,
fp32_1_A7,fp32_1_B7,
fp32_1_out
);

fp32PE fp32_2(clk,rst,
fp32_2_A0,fp32_2_B0,
fp32_2_A1,fp32_2_B1,
fp32_2_A2,fp32_2_B2,
fp32_2_A3,fp32_2_B3,
fp32_2_A4,fp32_2_B4,
fp32_2_A5,fp32_2_B5,
fp32_2_A6,fp32_2_B6,
fp32_2_A7,fp32_2_B7,
fp32_2_out
);

int8PE int8_0(clk,rst,
int8_0_A0,int8_0_B0,
int8_0_A1,int8_0_B1,
int8_0_A2,int8_0_B2,
int8_0_A3,int8_0_B3,
int8_0_A4,int8_0_B4,
int8_0_A5,int8_0_B5,
int8_0_A6,int8_0_B6,
int8_0_A7,int8_0_B7,
int8_0_out
);

int8PE int8_1(clk,rst,
int8_1_A0,int8_1_B0,
int8_1_A1,int8_1_B1,
int8_1_A2,int8_1_B2,
int8_1_A3,int8_1_B3,
int8_1_A4,int8_1_B4,
int8_1_A5,int8_1_B5,
int8_1_A6,int8_1_B6,
int8_1_A7,int8_1_B7,
int8_1_out
);

int8PE int8_2(clk,rst,
int8_2_A0,int8_2_B0,
int8_2_A1,int8_2_B1,
int8_2_A2,int8_2_B2,
int8_2_A3,int8_2_B3,
int8_2_A4,int8_2_B4,
int8_2_A5,int8_2_B5,
int8_2_A6,int8_2_B6,
int8_2_A7,int8_2_B7,
int8_2_out
);

mulPE muls0(
clk,
mulPE_0_ctrl,
mulPE_0_scalar,
mulPE_0_A0,mulPE_0_B0,
mulPE_0_A1,mulPE_0_B1,
mulPE_0_A2,mulPE_0_B2,
mulPE_0_A3,mulPE_0_B3,
mulPE_0_A4,mulPE_0_B4,
mulPE_0_A5,mulPE_0_B5,
mulPE_0_A6,mulPE_0_B6,
mulPE_0_A7,mulPE_0_B7,
mulPE_0_out0,
mulPE_0_out1,
mulPE_0_out2,
mulPE_0_out3,
mulPE_0_out4,
mulPE_0_out5,
mulPE_0_out6,
mulPE_0_out7
);

mulPE muls1(
clk,
mulPE_1_ctrl,
mulPE_1_scalar,
mulPE_1_A0,mulPE_1_B0,
mulPE_1_A1,mulPE_1_B1,
mulPE_1_A2,mulPE_1_B2,
mulPE_1_A3,mulPE_1_B3,
mulPE_1_A4,mulPE_1_B4,
mulPE_1_A5,mulPE_1_B5,
mulPE_1_A6,mulPE_1_B6,
mulPE_1_A7,mulPE_1_B7,
mulPE_1_out0,
mulPE_1_out1,
mulPE_1_out2,
mulPE_1_out3,
mulPE_1_out4,
mulPE_1_out5,
mulPE_1_out6,
mulPE_1_out7
);

mulPE muls2(
clk,
mulPE_2_ctrl,
mulPE_2_scalar,
mulPE_2_A0,mulPE_2_B0,
mulPE_2_A1,mulPE_2_B1,
mulPE_2_A2,mulPE_2_B2,
mulPE_2_A3,mulPE_2_B3,
mulPE_2_A4,mulPE_2_B4,
mulPE_2_A5,mulPE_2_B5,
mulPE_2_A6,mulPE_2_B6,
mulPE_2_A7,mulPE_2_B7,
mulPE_2_out0,
mulPE_2_out1,
mulPE_2_out2,
mulPE_2_out3,
mulPE_2_out4,
mulPE_2_out5,
mulPE_2_out6,
mulPE_2_out7
);

addPE adds0(
clk,
addPE_0_ctrl,
addPE_0_scalar,
addPE_0_A0,addPE_0_B0,
addPE_0_A1,addPE_0_B1,
addPE_0_A2,addPE_0_B2,
addPE_0_A3,addPE_0_B3,
addPE_0_A4,addPE_0_B4,
addPE_0_A5,addPE_0_B5,
addPE_0_A6,addPE_0_B6,
addPE_0_A7,addPE_0_B7,
addPE_0_out0,
addPE_0_out1,
addPE_0_out2,
addPE_0_out3,
addPE_0_out4,
addPE_0_out5,
addPE_0_out6,
addPE_0_out7
);

addPE adds1(
clk,
addPE_1_ctrl,
addPE_1_scalar,
addPE_1_A0,addPE_1_B0,
addPE_1_A1,addPE_1_B1,
addPE_1_A2,addPE_1_B2,
addPE_1_A3,addPE_1_B3,
addPE_1_A4,addPE_1_B4,
addPE_1_A5,addPE_1_B5,
addPE_1_A6,addPE_1_B6,
addPE_1_A7,addPE_1_B7,
addPE_1_out0,
addPE_1_out1,
addPE_1_out2,
addPE_1_out3,
addPE_1_out4,
addPE_1_out5,
addPE_1_out6,
addPE_1_out7
);

addPE adds2(
clk,
addPE_2_ctrl,
addPE_2_scalar,
addPE_2_A0,addPE_2_B0,
addPE_2_A1,addPE_2_B1,
addPE_2_A2,addPE_2_B2,
addPE_2_A3,addPE_2_B3,
addPE_2_A4,addPE_2_B4,
addPE_2_A5,addPE_2_B5,
addPE_2_A6,addPE_2_B6,
addPE_2_A7,addPE_2_B7,
addPE_2_out0,
addPE_2_out1,
addPE_2_out2,
addPE_2_out3,
addPE_2_out4,
addPE_2_out5,
addPE_2_out6,
addPE_2_out7
);

treePE trees0(
clk,
rst,
treePE_0_A0,
treePE_0_A1,
treePE_0_A2,
treePE_0_A3,
treePE_0_A4,
treePE_0_A5,
treePE_0_A6,
treePE_0_A7,
treePE_0_out
);

treePE trees1(
clk,
rst,
treePE_1_A0,
treePE_1_A1,
treePE_1_A2,
treePE_1_A3,
treePE_1_A4,
treePE_1_A5,
treePE_1_A6,
treePE_1_A7,
treePE_1_out
);

treePE trees2(
clk,
rst,
treePE_2_A0,
treePE_2_A1,
treePE_2_A2,
treePE_2_A3,
treePE_2_A4,
treePE_2_A5,
treePE_2_A6,
treePE_2_A7,
treePE_2_out
);

endmodule